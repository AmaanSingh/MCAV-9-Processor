//go from instr_rom to decoder to control and reg file