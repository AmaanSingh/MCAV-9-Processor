//go from instr_rom to decoder to control and reg file
module decoder (
  input					clk,
  input					rst,
  input					instruction_decode_en,

  // to register file
  output          [7:0] dat_in,
  
);  



endmodule